module test_temp #(parameter aa=1) (
  input clk, //input clk
  input rst_n,
  output [31:0] data_in,
  input done
);

wire test;
wire test1;

assign test = test1;

endmodule

