module test_temp_1 #(parameter aa=1) (
  input rst_n,
  input [31:0] data_in,
  output [31:0] data_out,
  output done
);

wire test;
wire test1;

assign test = test1;

endmodule

