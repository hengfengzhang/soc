module test_temp #(parameter aa=1) (
  input clk, //input clk
  input rst_n,
  input [31:0] data_in,
  output done
);

wire test;
wire test1;

assign test = test1;

endmodule

